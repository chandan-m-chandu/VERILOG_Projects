module full_adder(input wire A,B,Cin, output wire Y);
  assign Y = A^B^Cin;
endmodule
